// ===========================================================================
// Restricted (c) Siemens 2024. 
// All Rights Reserved 
// THIS WORK CONTAINS TRADE SECRET AND CONFIDENTIAL INFORMATION WHICH ARE THE PROPERTY OF 
// MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO LICENSE TERMS. 
//
// File description: Evaluation subsystem.
//
// Customer modification rights are granted for this file.
//
// ===========================================================================

`include "ust_defines.vh"
//`include "ust_std.vh"
module ust_ss_bosc_eval_m
  #(
  parameter index_length_p = 8,
  parameter me0_clk_disable_reset_p = 1,
  parameter me0_gpio_in_width_p = 8,
  parameter me0_gpio_out_width_p = 8,
  parameter me0_gpio_p = 0,
  parameter me0_gpio_reset_p = 0,
  parameter me0_hysteresis_width_p = 0,
  parameter me0_info_width_p = 8,
  parameter me0_pipeline_p = 0,
  parameter me0_time_p = 1,
  parameter me0_lower_0_bypass_p = 1,
  parameter me0_lower_0_ingress_event_depth_p = 1,
  parameter me0_lower_0_ingress_msg_depth_p = 0,
  parameter me0_lower_0_egress_msg_depth_p = 0,
  parameter me0_lower_0_event_mask_width_p = 0,
  parameter me0_upper_0_bypass_p = 1,
  parameter me0_upper_0_ingress_event_depth_p = 1,
  parameter me0_upper_0_ingress_msg_depth_p = 0,
  parameter me0_upper_0_egress_msg_depth_p = 0,
  parameter me0_upper_0_event_mask_width_p = 0,
  parameter me0_upper_1_bypass_p = 1,
  parameter me0_upper_1_ingress_event_depth_p = 1,
  parameter me0_upper_1_ingress_msg_depth_p = 0,
  parameter me0_upper_1_egress_msg_depth_p = 0,
  parameter me0_upper_1_event_mask_width_p = 0,
  parameter lower_0_us_msg_sz_p = 5,
  parameter lower_0_ds_msg_sz_p = 5,
  parameter ete0_auth_p = 0,
  parameter ete0_alloc_p = 0,
  parameter ete0_bypass_p = 0,
  parameter ete0_comparators_p = 2,
  parameter ete0_counters_p = 0,
  parameter ete0_counter_width_p = 16,
  parameter ete0_filters_p = 1,
  parameter ete0_trace_bypass_p = 0,
  parameter ete0_itrace_size_p = 128,
  parameter ete0_itrace_fast_p = 0,
  parameter ete0_lossless_p = 0,
  parameter ete0_nocontext_p = 1,
  parameter ete0_context_width_p = 32,
  parameter ete0_ctype_width_p = 2,
  parameter ete0_ecause_width_p = 5,
  parameter ete0_ecause_choice_p = 5,
  parameter ete0_impexcept_p = 2,
  parameter ete0_iaddress_lsb_p = 1,
  parameter ete0_iaddress_width_p = 32,
  parameter ete0_lastsize_linear_p = 0,
  parameter ete0_lastsize_width_p = 1,
  parameter ete0_nodiffaddr_p = 0,
  parameter ete0_itype_width_p = 4,
  parameter ete0_privilege_width_p = 2,
  parameter ete0_privilege_reset_p = 3,
  parameter ete0_sijump_p = 0,
  parameter ete0_uiret_p = 0,
  parameter ete0_bpred_size_p = 0,
  parameter ete0_cache_size_p = 0,
  parameter ete0_call_counter_size_p = 0,
  parameter ete0_return_stack_size_p = 0,
  parameter ete0_status_width_p = 1,
  parameter ete0_impdef_width_p = 1,
  parameter ete0_filter_iaddress_p = 1,
  parameter ete0_filter_context_p = 1,
  parameter ete0_filter_excint_p = 1,
  parameter ete0_filter_privilege_p = 1,
  parameter ete0_filter_tval_p = 1,
  parameter ete0_filter_impdef_p = 1,
  parameter ete0_ds_msg_sz_p = 5,
  parameter ete0_us_msg_sz_p = 3,
  parameter ete0_us_cdc_depth_p = 0,
  parameter ete0_ds_event_fifo_depth_p = 4,
  parameter ete0_pipeline_p = 1,
  parameter ete0_timer_width_p = 32,
  parameter ete0_gpio_p = 1,
  parameter ete0_gpio_out_width_p = 8,
  parameter ete0_gpio_reset_p = 0,
  parameter ete0_test_0_mtype_p = 1,
  parameter ete0_test_in_0_width_p = 1,
  parameter ete0_test_out_0_width_p = 1,
  parameter ete0_udb2sys_sync_stages_p = 2,
  parameter ete0_sys2udb_sync_stages_p = 2,
  parameter ust_upper_0_indexes_p = 1,
  parameter ete_mult_retire_auth_p = 0,
  parameter ete_mult_retire_alloc_p = 0,
  parameter ete_mult_retire_bypass_p = 1,
  parameter ete_mult_retire_comparators_p = 2,
  parameter ete_mult_retire_counters_p = 0,
  parameter ete_mult_retire_counter_width_p = 16,
  parameter ete_mult_retire_filters_p = 1,
  parameter ete_mult_retire_trace_bypass_p = 1,
  parameter ete_mult_retire_itrace_size_p = 128,
  parameter ete_mult_retire_itrace_fast_p = 0,
  parameter ete_mult_retire_lossless_p = 0,
  parameter ete_mult_retire_nocontext_p = 0,
  parameter ete_mult_retire_context_width_p = 32,
  parameter ete_mult_retire_ctype_width_p = 2,
  parameter ete_mult_retire_ecause_width_p = 5,
  parameter ete_mult_retire_ecause_choice_p = 5,
  parameter ete_mult_retire_impexcept_p = 2,
  parameter ete_mult_retire_iaddress_lsb_p = 1,
  parameter ete_mult_retire_iaddress_width_p = 32,
  parameter ete_mult_retire_lastsize_linear_p = 0,
  parameter ete_mult_retire_lastsize_width_p = 1,
  parameter ete_mult_retire_nodiffaddr_p = 0,
  parameter ete_mult_retire_itype_width_p = 4,
  parameter ete_mult_retire_privilege_width_p = 4,
  parameter ete_mult_retire_privilege_reset_p = 0,
  parameter ete_mult_retire_sijump_p = 1,
  parameter ete_mult_retire_uiret_p = 0,
  parameter ete_mult_retire_bpred_size_p = 0,
  parameter ete_mult_retire_cache_size_p = 0,
  parameter ete_mult_retire_call_counter_size_p = 0,
  parameter ete_mult_retire_return_stack_size_p = 0,
  parameter ete_mult_retire_status_width_p = 4,
  parameter ete_mult_retire_impdef_width_p = 1,
  parameter ete_mult_retire_filter_iaddress_p = 1,
  parameter ete_mult_retire_filter_context_p = 1,
  parameter ete_mult_retire_filter_excint_p = 1,
  parameter ete_mult_retire_filter_privilege_p = 1,
  parameter ete_mult_retire_filter_tval_p = 1,
  parameter ete_mult_retire_filter_impdef_p = 1,
  parameter ete_mult_retire_ds_msg_sz_p = 5,
  parameter ete_mult_retire_us_msg_sz_p = 3,
  parameter ete_mult_retire_us_cdc_depth_p = 0,
  parameter ete_mult_retire_ds_event_fifo_depth_p = 4,
  parameter ete_mult_retire_pipeline_p = 0,
  parameter ete_mult_retire_timer_width_p = 32,
  parameter ete_mult_retire_gpio_p = 1,
  parameter ete_mult_retire_gpio_out_width_p = 8,
  parameter ete_mult_retire_gpio_reset_p = 0,
  parameter ete_mult_retire_test_0_mtype_p = 1,
  parameter ete_mult_retire_test_in_0_width_p = 1,
  parameter ete_mult_retire_test_out_0_width_p = 1,
  parameter ete_mult_retire_udb2sys_sync_stages_p = 2,
  parameter ete_mult_retire_sys2udb_sync_stages_p = 2,
  parameter ete_mult_retire_iblocks_p = 1,
  parameter ete_mult_retire_iretires_p = 2,
  parameter ust_upper_1_indexes_p = 1,
  parameter ete0_iretires_p = 1
  )
  (
  input wire   ust_clk_udb_ip,
  input wire   ust_rst_udb_ip,
  output wire [(me0_gpio_out_width_p)-1:0] ust_me0_gpio_out_op,
  input  wire [(me0_gpio_in_width_p)-1:0]  ust_me0_gpio_in_ip,
  input wire [15:0] ust_me0_instance_id_ip,
  input wire [31:0] ust_me0_idcode_ip,
  input wire [(index_length_p)-1:0] ust_me0_msg_reserved_ip,
  input wire [(me0_info_width_p)-1:0] ust_me0_chip_info_ip,
  output wire [31:0] ust_me0_time_op,
  input wire [3:0] ust_me0_flow0_route_ip,
  input wire [3:0] ust_me0_flow1_route_ip,
  input wire [3:0] ust_me0_flow2_route_ip,
  input  wire [(2**lower_0_us_msg_sz_p)-1:0] ust_lower_0_us_msg_data_ip,
  input  wire                                ust_lower_0_us_msg_event_ip,
  output wire                                ust_lower_0_us_msg_ready_op,
  input  wire                                ust_lower_0_us_msg_valid_ip,
  output wire [(2**lower_0_ds_msg_sz_p)-1:0] ust_lower_0_ds_msg_data_op,
  output wire                                ust_lower_0_ds_msg_event_op,
  input  wire                                ust_lower_0_ds_msg_ready_ip,
  output wire                                ust_lower_0_ds_msg_valid_op,
  input  wire                                ust_ete0_rv_halted_ip,// Halted
  output wire                                ust_ete0_rv_stall_op,  // Stall
  input  wire [(1)-1:0]                      ust_ete0_rv_i_retire_ip,// Number of halfwords retired
  input  wire [(ete0_lastsize_width_p)-1:0]  ust_ete0_rv_i_lastsize_ip,// Size of last instruction in block is 2**ust_rv_i_lastsize_ip halfwords
  input  wire [(ete0_itype_width_p)-1:0]     ust_ete0_rv_i_type_ip,  // Type of last retired instruction
  input  wire [(1)-1:0]                      ust_ete0_rv_i_sijump_ip,// Last retired instruction is a sequentially inferable jump
  input  wire [(ete0_iaddress_width_p)-1:0]  ust_ete0_rv_i_address_ip,// Instruction address
  input  wire [(ete0_context_width_p)-1:0]   ust_ete0_rv_i_context_ip,// Instruction context
  input  wire [(ete0_ctype_width_p)-1:0]     ust_ete0_rv_i_ctype_ip,// Instruction context type
  input  wire [(ete0_ecause_width_p)-1:0]    ust_ete0_rv_i_ecause_ip,// Exception cause
  input  wire [(ete0_iaddress_width_p)-1:0]  ust_ete0_rv_i_tval_ip,// Exception trap value
  input  wire [(ete0_privilege_width_p)-1:0] ust_ete0_rv_i_privilege_ip,// Privilege level
  input  wire [(3)-1:0]                      ust_ete0_rv_i_trigger_ip,// Debug Module triggers (bit 2 replicated per block)
  input  wire [(ete0_impdef_width_p)-1:0]    ust_ete0_rv_i_impdef_ip,// Implementation-defined filter qualifiers
  input  wire [(ete0_status_width_p)-1:0]    ust_ete0_rv_i_status_ip,
  output wire                                ust_ete0_rv_i_enabled_op,// Enabled
  input wire   ust_clk_ete0_sys_ip,
  input wire   ust_rst_ete0_sys_ip,
  output wire   ust_en_ete0_sys_op,
  input wire   ust_ete0_testmode_ip,
  output wire [(ete0_gpio_out_width_p)-1:0] ust_ete0_gpio_output_op,
  output wire [8:0] ust_ete0_version_op,
  input wire [15:0] ust_ete0_instance_id_ip,
  input  wire                                                                                                                                                   ust_ete_mult_retire_rv_halted_ip,     // Halted
  output wire                                                                                                                                                   ust_ete_mult_retire_rv_stall_op,// Stall
  input  wire [(ete_mult_retire_iretires_p > 1 ? ete_mult_retire_iblocks_p * `ust_clog2((ete_mult_retire_iretires_p * 2) + 1) : ete_mult_retire_iblocks_p)-1:0] ust_ete_mult_retire_rv_i_retire_ip,  //Number of halfwords retired
  input  wire [(ete_mult_retire_iblocks_p * ete_mult_retire_lastsize_width_p)-1:0]                                                                              ust_ete_mult_retire_rv_i_lastsize_ip,//Size of last instruction in block is 2**ust_rv_i_lastsize_ip halfwords
  input  wire [(ete_mult_retire_iblocks_p * ete_mult_retire_itype_width_p)-1:0]                                                                                 ust_ete_mult_retire_rv_i_type_ip, // Type of last retired instruction
  input  wire [(ete_mult_retire_iblocks_p)-1:0]                                                                                                                 ust_ete_mult_retire_rv_i_sijump_ip,// Last retired instruction is a sequentially inferable jump
  input  wire [(ete_mult_retire_iblocks_p)-1:0]                                                                                                                 ust_ete_mult_retire_rv_i_uiret_ip,
  input  wire [(ete_mult_retire_iblocks_p * ete_mult_retire_iaddress_width_p)-1:0]                                                                              ust_ete_mult_retire_rv_i_address_ip,// Instruction address
  input  wire [(ete_mult_retire_context_width_p)-1:0]                                                                                                           ust_ete_mult_retire_rv_i_context_ip,// Instruction context type
  input  wire [(ete_mult_retire_ctype_width_p)-1:0]                                                                                                             ust_ete_mult_retire_rv_i_ctype_ip,
  input  wire [(ete_mult_retire_ecause_width_p)-1:0]                                                                                                            ust_ete_mult_retire_rv_i_ecause_ip,// Exception cause
  input  wire [(ete_mult_retire_iaddress_width_p)-1:0]                                                                                                          ust_ete_mult_retire_rv_i_tval_ip,// Exception trap value
  input  wire [(ete_mult_retire_privilege_width_p)-1:0]                                                                                                         ust_ete_mult_retire_rv_i_privilege_ip,// Privilege level
  input  wire [(2 + ete_mult_retire_iblocks_p)-1:0]                                                                                                             ust_ete_mult_retire_rv_i_trigger_ip,// Debug Module triggers (bit 2 replicated per block)
  input  wire [(ete_mult_retire_impdef_width_p)-1:0]                                                                                                            ust_ete_mult_retire_rv_i_impdef_ip,// Implementation-defined filter qualifiers
  input  wire [(ete_mult_retire_status_width_p)-1:0]                                                                                                            ust_ete_mult_retire_rv_i_status_ip,// Status flags
  output wire                                                                                                                                                   ust_ete_mult_retire_rv_i_enabled_op,// Enabled
  input wire   ust_clk_ete_mult_retire_sys_ip,
  input wire   ust_rst_ete_mult_retire_sys_ip,
  output wire   ust_en_ete_mult_retire_sys_op,
  input wire   ust_ete_mult_retire_testmode_ip,
  output wire [(ete_mult_retire_gpio_out_width_p)-1:0] ust_ete_mult_retire_gpio_output_op,
  output wire [8:0] ust_ete_mult_retire_version_op,
  input wire [15:0] ust_ete_mult_retire_instance_id_ip
  );
  
  
  wire [(1)-1:0] _dummy_w;
  
  wire [(2**ete0_us_msg_sz_p)-1:0] ust_ete0_us_msg_data_w;
  wire                             ust_ete0_us_msg_event_w;
  wire                             ust_ete0_us_msg_ready_w;
  wire                             ust_ete0_us_msg_valid_w;
  wire [(2**ete0_ds_msg_sz_p)-1:0] ust_ete0_ds_msg_data_w;
  wire                             ust_ete0_ds_msg_event_w;
  wire                             ust_ete0_ds_msg_ready_w;
  wire                             ust_ete0_ds_msg_valid_w;
  
  wire [(2**ete_mult_retire_us_msg_sz_p)-1:0] ust_ete_mult_retire_us_msg_data_w;
  wire                                        ust_ete_mult_retire_us_msg_event_w;
  wire                                        ust_ete_mult_retire_us_msg_ready_w;
  wire                                        ust_ete_mult_retire_us_msg_valid_w;
  wire [(2**ete_mult_retire_ds_msg_sz_p)-1:0] ust_ete_mult_retire_ds_msg_data_w;
  wire                                        ust_ete_mult_retire_ds_msg_event_w;
  wire                                        ust_ete_mult_retire_ds_msg_ready_w;
  wire                                        ust_ete_mult_retire_ds_msg_valid_w;
  
  ust_me_l1u2s0_m
   #(
    .index_length_p                ( index_length_p                    ),
    .clk_disable_reset_p           ( me0_clk_disable_reset_p           ),
    .cm_support_p                  ( 0                                 ),
    .gpio_in_width_p               ( me0_gpio_in_width_p               ),
    .gpio_out_width_p              ( me0_gpio_out_width_p              ),
    .gpio_p                        ( me0_gpio_p                        ),
    .gpio_reset_p                  ( me0_gpio_reset_p                  ),
    .hysteresis_width_p            ( me0_hysteresis_width_p            ),
    .info_width_p                  ( me0_info_width_p                  ),
    .pipeline_p                    ( me0_pipeline_p                    ),
    .time_p                        ( me0_time_p                        ),
    .lower_0_bypass_p              ( me0_lower_0_bypass_p              ),
    .lower_0_ds_msg_sz_p           ( lower_0_ds_msg_sz_p               ),
    .lower_0_us_msg_sz_p           ( lower_0_us_msg_sz_p               ),
    .lower_0_ingress_event_depth_p ( me0_lower_0_ingress_event_depth_p ),
    .lower_0_ingress_msg_depth_p   ( me0_lower_0_ingress_msg_depth_p   ),
    .lower_0_egress_msg_depth_p    ( me0_lower_0_egress_msg_depth_p    ),
    .lower_0_event_mask_width_p    ( me0_lower_0_event_mask_width_p    ),
    .upper_0_bypass_p              ( me0_upper_0_bypass_p              ),
    .upper_0_ds_msg_sz_p           ( ete0_ds_msg_sz_p                  ),
    .upper_0_us_msg_sz_p           ( ete0_us_msg_sz_p                  ),
    .upper_0_ingress_event_depth_p ( me0_upper_0_ingress_event_depth_p ),
    .upper_0_ingress_msg_depth_p   ( me0_upper_0_ingress_msg_depth_p   ),
    .upper_0_egress_msg_depth_p    ( me0_upper_0_egress_msg_depth_p    ),
    .upper_0_event_mask_width_p    ( me0_upper_0_event_mask_width_p    ),
    .upper_1_bypass_p              ( me0_upper_1_bypass_p              ),
    .upper_1_ds_msg_sz_p           ( ete_mult_retire_ds_msg_sz_p       ),
    .upper_1_us_msg_sz_p           ( ete_mult_retire_us_msg_sz_p       ),
    .upper_1_ingress_event_depth_p ( me0_upper_1_ingress_event_depth_p ),
    .upper_1_ingress_msg_depth_p   ( me0_upper_1_ingress_msg_depth_p   ),
    .upper_1_egress_msg_depth_p    ( me0_upper_1_egress_msg_depth_p    ),
    .upper_1_event_mask_width_p    ( me0_upper_1_event_mask_width_p    )
  ) 
  me0 (
    .ust_clk_udb_ip              ( ust_clk_udb_ip                             ),
    .ust_rst_udb_ip              ( ust_rst_udb_ip                             ),
    .ust_instance_id_ip          ( ust_me0_instance_id_ip                     ),
    .ust_idcode_ip               ( ust_me0_idcode_ip                          ),
    .ust_chip_info_ip            ( ust_me0_chip_info_ip                       ),
    .ust_msg_reserved_ip         ( ust_me0_msg_reserved_ip                    ),
    .ust_time_op                 ( ust_me0_time_op                            ),
    .ust_gpio_out_op             ( ust_me0_gpio_out_op                        ),
    .ust_gpio_in_ip              ( ust_me0_gpio_in_ip                         ),
    .ust_msg_indexes_op          (                                            ),
    .ust_flow0_route_ip          ( ust_me0_flow0_route_ip                     ),
    .ust_flow1_route_ip          ( ust_me0_flow1_route_ip                     ),
    .ust_flow2_route_ip          ( ust_me0_flow2_route_ip                     ),
    .ust_lower_0_indexes_ip      ( {(index_length_p){1'b0}}                   ),
    .ust_lower_0_us_msg_data_ip  ( ust_lower_0_us_msg_data_ip                 ),
    .ust_lower_0_us_msg_event_ip ( ust_lower_0_us_msg_event_ip                ),
    .ust_lower_0_us_msg_ready_op ( ust_lower_0_us_msg_ready_op                ),
    .ust_lower_0_us_msg_valid_ip ( ust_lower_0_us_msg_valid_ip                ),
    .ust_lower_0_ds_msg_data_op  ( ust_lower_0_ds_msg_data_op                 ),
    .ust_lower_0_ds_msg_event_op ( ust_lower_0_ds_msg_event_op                ),
    .ust_lower_0_ds_msg_ready_ip ( ust_lower_0_ds_msg_ready_ip                ),
    .ust_lower_0_ds_msg_valid_op ( ust_lower_0_ds_msg_valid_op                ),
    .ust_upper_0_indexes_ip      ( ust_upper_0_indexes_p[index_length_p-1:0]  ),
    .ust_upper_0_us_msg_data_op  ( ust_ete0_us_msg_data_w                     ),
    .ust_upper_0_us_msg_event_op ( ust_ete0_us_msg_event_w                    ),
    .ust_upper_0_us_msg_ready_ip ( ust_ete0_us_msg_ready_w                    ),
    .ust_upper_0_us_msg_valid_op ( ust_ete0_us_msg_valid_w                    ),
    .ust_upper_0_ds_msg_data_ip  ( ust_ete0_ds_msg_data_w                     ),
    .ust_upper_0_ds_msg_event_ip ( ust_ete0_ds_msg_event_w                    ),
    .ust_upper_0_ds_msg_ready_op ( ust_ete0_ds_msg_ready_w                    ),
    .ust_upper_0_ds_msg_valid_ip ( ust_ete0_ds_msg_valid_w                    ),
    .ust_upper_1_indexes_ip      ( ust_upper_1_indexes_p[index_length_p-1:0]  ),
    .ust_upper_1_us_msg_data_op  ( ust_ete_mult_retire_us_msg_data_w          ),
    .ust_upper_1_us_msg_event_op ( ust_ete_mult_retire_us_msg_event_w         ),
    .ust_upper_1_us_msg_ready_ip ( ust_ete_mult_retire_us_msg_ready_w         ),
    .ust_upper_1_us_msg_valid_op ( ust_ete_mult_retire_us_msg_valid_w         ),
    .ust_upper_1_ds_msg_data_ip  ( ust_ete_mult_retire_ds_msg_data_w          ),
    .ust_upper_1_ds_msg_event_ip ( ust_ete_mult_retire_ds_msg_event_w         ),
    .ust_upper_1_ds_msg_ready_op ( ust_ete_mult_retire_ds_msg_ready_w         ),
    .ust_upper_1_ds_msg_valid_ip ( ust_ete_mult_retire_ds_msg_valid_w         )
  );
  
  
  ust_etrace_encoder_a0t1_m
   #(
    .index_length_p        ( index_length_p             ),
    .auth_p                ( ete0_auth_p                ),
    .alloc_p               ( ete0_alloc_p               ),
    .bypass_p              ( ete0_bypass_p              ),
    .comparators_p         ( ete0_comparators_p         ),
    .counters_p            ( ete0_counters_p            ),
    .counter_width_p       ( ete0_counter_width_p       ),
    .filters_p             ( ete0_filters_p             ),
    .trace_bypass_p        ( ete0_trace_bypass_p        ),
    .itrace_size_p         ( ete0_itrace_size_p         ),
    .itrace_fast_p         ( ete0_itrace_fast_p         ),
    .lossless_p            ( ete0_lossless_p            ),
    .nocontext_p           ( ete0_nocontext_p           ),
    .context_width_p       ( ete0_context_width_p       ),
    .ctype_width_p         ( ete0_ctype_width_p         ),
    .ecause_width_p        ( ete0_ecause_width_p        ),
    .ecause_choice_p       ( ete0_ecause_choice_p       ),
    .impexcept_p           ( ete0_impexcept_p           ),
    .iaddress_lsb_p        ( ete0_iaddress_lsb_p        ),
    .iaddress_width_p      ( ete0_iaddress_width_p      ),
    .lastsize_linear_p     ( ete0_lastsize_linear_p     ),
    .lastsize_width_p      ( ete0_lastsize_width_p      ),
    .nodiffaddr_p          ( ete0_nodiffaddr_p          ),
    .itype_width_p         ( ete0_itype_width_p         ),
    .privilege_width_p     ( ete0_privilege_width_p     ),
    .privilege_reset_p     ( ete0_privilege_reset_p     ),
    .sijump_p              ( ete0_sijump_p              ),
    .uiret_p               ( ete0_uiret_p               ),
    .bpred_size_p          ( ete0_bpred_size_p          ),
    .cache_size_p          ( ete0_cache_size_p          ),
    .call_counter_size_p   ( ete0_call_counter_size_p   ),
    .return_stack_size_p   ( ete0_return_stack_size_p   ),
    .status_width_p        ( ete0_status_width_p        ),
    .impdef_width_p        ( ete0_impdef_width_p        ),
    .filter_iaddress_p     ( ete0_filter_iaddress_p     ),
    .filter_context_p      ( ete0_filter_context_p      ),
    .filter_excint_p       ( ete0_filter_excint_p       ),
    .filter_privilege_p    ( ete0_filter_privilege_p    ),
    .filter_tval_p         ( ete0_filter_tval_p         ),
    .filter_impdef_p       ( ete0_filter_impdef_p       ),
    .ds_msg_sz_p           ( ete0_ds_msg_sz_p           ),
    .us_msg_sz_p           ( ete0_us_msg_sz_p           ),
    .us_cdc_depth_p        ( ete0_us_cdc_depth_p        ),
    .ds_event_fifo_depth_p ( ete0_ds_event_fifo_depth_p ),
    .pipeline_p            ( ete0_pipeline_p            ),
    .timer_width_p         ( ete0_timer_width_p         ),
    .gpio_p                ( ete0_gpio_p                ),
    .gpio_out_width_p      ( ete0_gpio_out_width_p      ),
    .gpio_reset_p          ( ete0_gpio_reset_p          ),
    .test_0_mtype_p        ( ete0_test_0_mtype_p        ),
    .test_in_0_width_p     ( ete0_test_in_0_width_p     ),
    .test_out_0_width_p    ( ete0_test_out_0_width_p    ),
    .udb2sys_sync_stages_p ( ete0_udb2sys_sync_stages_p ),
    .sys2udb_sync_stages_p ( ete0_sys2udb_sync_stages_p )
  ) 
  ete0 (
    .ust_clk_udb_ip        ( ust_clk_udb_ip                    ),
    .ust_rst_udb_ip        ( ust_rst_udb_ip                    ),
    .ust_clk_sys_ip        ( ust_clk_ete0_sys_ip               ),
    .ust_rst_sys_ip        ( ust_rst_ete0_sys_ip               ),
    .ust_en_sys_op         ( ust_en_ete0_sys_op                ),
    .ust_us_msg_data_ip    ( ust_ete0_us_msg_data_w            ),
    .ust_us_msg_event_ip   ( ust_ete0_us_msg_event_w           ),
    .ust_us_msg_ready_op   ( ust_ete0_us_msg_ready_w           ),
    .ust_us_msg_valid_ip   ( ust_ete0_us_msg_valid_w           ),
    .ust_ds_msg_data_op    ( ust_ete0_ds_msg_data_w            ),
    .ust_ds_msg_event_op   ( ust_ete0_ds_msg_event_w           ),
    .ust_ds_msg_ready_ip   ( ust_ete0_ds_msg_ready_w           ),
    .ust_ds_msg_valid_op   ( ust_ete0_ds_msg_valid_w           ),
    .ust_gpio_output_op    ( ust_ete0_gpio_output_op           ),
    .ust_rv_halted_ip      ( ust_ete0_rv_halted_ip             ),
    .ust_rv_stall_op       ( ust_ete0_rv_stall_op              ),
    .ust_rv_i_retire_ip    ( ust_ete0_rv_i_retire_ip           ),
    .ust_rv_i_lastsize_ip  ( ust_ete0_rv_i_lastsize_ip         ),
    .ust_rv_i_type_ip      ( ust_ete0_rv_i_type_ip             ),
    .ust_rv_i_sijump_ip    ( ust_ete0_rv_i_sijump_ip           ),
    .ust_rv_i_uiret_ip     ( ust_ete0_rv_i_uiret_ip            ),
    .ust_rv_i_address_ip   ( ust_ete0_rv_i_address_ip          ),
    .ust_rv_i_context_ip   ( ust_ete0_rv_i_context_ip          ),
    .ust_rv_i_ctype_ip     ( ust_ete0_rv_i_ctype_ip            ),
    .ust_rv_i_ecause_ip    ( ust_ete0_rv_i_ecause_ip           ),
    .ust_rv_i_tval_ip      ( ust_ete0_rv_i_tval_ip             ),
    .ust_rv_i_privilege_ip ( ust_ete0_rv_i_privilege_ip        ),
    .ust_rv_i_trigger_ip   ( ust_ete0_rv_i_trigger_ip          ),
    .ust_rv_i_impdef_ip    ( ust_ete0_rv_i_impdef_ip           ),
    .ust_rv_i_status_ip    ( ust_ete0_rv_i_status_ip           ),
    .ust_rv_i_enabled_op   ( ust_ete0_rv_i_enabled_op          ),
    .ust_lock_ip           ( 1'd0                              ),
    .ust_locked_op         (                                   ),
    .ust_instance_id_ip    ( ust_ete0_instance_id_ip           ),
    .ust_version_op        ( ust_ete0_version_op               ),
    .ust_testmode_ip       ( ust_ete0_testmode_ip              ),
    .ust_test_in_0_ip      ( {(ete0_test_in_0_width_p){1'b0}}  ),
    .ust_test_out_0_op     (                                   )
  );
  
  ust_etrace_encoder_a1t1_m
   #(
    .index_length_p        ( index_length_p                        ),
    .auth_p                ( ete_mult_retire_auth_p                ),
    .alloc_p               ( ete_mult_retire_alloc_p               ),
    .bypass_p              ( ete_mult_retire_bypass_p              ),
    .comparators_p         ( ete_mult_retire_comparators_p         ),
    .counters_p            ( ete_mult_retire_counters_p            ),
    .counter_width_p       ( ete_mult_retire_counter_width_p       ),
    .filters_p             ( ete_mult_retire_filters_p             ),
    .trace_bypass_p        ( ete_mult_retire_trace_bypass_p        ),
    .itrace_size_p         ( ete_mult_retire_itrace_size_p         ),
    .itrace_fast_p         ( ete_mult_retire_itrace_fast_p         ),
    .lossless_p            ( ete_mult_retire_lossless_p            ),
    .nocontext_p           ( ete_mult_retire_nocontext_p           ),
    .context_width_p       ( ete_mult_retire_context_width_p       ),
    .ctype_width_p         ( ete_mult_retire_ctype_width_p         ),
    .ecause_width_p        ( ete_mult_retire_ecause_width_p        ),
    .ecause_choice_p       ( ete_mult_retire_ecause_choice_p       ),
    .impexcept_p           ( ete_mult_retire_impexcept_p           ),
    .iaddress_lsb_p        ( ete_mult_retire_iaddress_lsb_p        ),
    .iaddress_width_p      ( ete_mult_retire_iaddress_width_p      ),
    .lastsize_linear_p     ( ete_mult_retire_lastsize_linear_p     ),
    .lastsize_width_p      ( ete_mult_retire_lastsize_width_p      ),
    .nodiffaddr_p          ( ete_mult_retire_nodiffaddr_p          ),
    .itype_width_p         ( ete_mult_retire_itype_width_p         ),
    .privilege_width_p     ( ete_mult_retire_privilege_width_p     ),
    .privilege_reset_p     ( ete_mult_retire_privilege_reset_p     ),
    .sijump_p              ( ete_mult_retire_sijump_p              ),
    .uiret_p               ( ete_mult_retire_uiret_p               ),
    .bpred_size_p          ( ete_mult_retire_bpred_size_p          ),
    .cache_size_p          ( ete_mult_retire_cache_size_p          ),
    .call_counter_size_p   ( ete_mult_retire_call_counter_size_p   ),
    .return_stack_size_p   ( ete_mult_retire_return_stack_size_p   ),
    .status_width_p        ( ete_mult_retire_status_width_p        ),
    .impdef_width_p        ( ete_mult_retire_impdef_width_p        ),
    .filter_iaddress_p     ( ete_mult_retire_filter_iaddress_p     ),
    .filter_context_p      ( ete_mult_retire_filter_context_p      ),
    .filter_excint_p       ( ete_mult_retire_filter_excint_p       ),
    .filter_privilege_p    ( ete_mult_retire_filter_privilege_p    ),
    .filter_tval_p         ( ete_mult_retire_filter_tval_p         ),
    .filter_impdef_p       ( ete_mult_retire_filter_impdef_p       ),
    .ds_msg_sz_p           ( ete_mult_retire_ds_msg_sz_p           ),
    .us_msg_sz_p           ( ete_mult_retire_us_msg_sz_p           ),
    .us_cdc_depth_p        ( ete_mult_retire_us_cdc_depth_p        ),
    .ds_event_fifo_depth_p ( ete_mult_retire_ds_event_fifo_depth_p ),
    .pipeline_p            ( ete_mult_retire_pipeline_p            ),
    .timer_width_p         ( ete_mult_retire_timer_width_p         ),
    .gpio_p                ( ete_mult_retire_gpio_p                ),
    .gpio_out_width_p      ( ete_mult_retire_gpio_out_width_p      ),
    .gpio_reset_p          ( ete_mult_retire_gpio_reset_p          ),
    .test_0_mtype_p        ( ete_mult_retire_test_0_mtype_p        ),
    .test_in_0_width_p     ( ete_mult_retire_test_in_0_width_p     ),
    .test_out_0_width_p    ( ete_mult_retire_test_out_0_width_p    ),
    .udb2sys_sync_stages_p ( ete_mult_retire_udb2sys_sync_stages_p ),
    .sys2udb_sync_stages_p ( ete_mult_retire_sys2udb_sync_stages_p ),
    .iblocks_p             ( ete_mult_retire_iblocks_p             ),
    .iretires_p            ( ete_mult_retire_iretires_p            )
  ) 
  ete_mult_retire (
    .ust_clk_udb_ip        ( ust_clk_udb_ip                               ),
    .ust_rst_udb_ip        ( ust_rst_udb_ip                               ),
    .ust_clk_sys_ip        ( ust_clk_ete_mult_retire_sys_ip               ),
    .ust_rst_sys_ip        ( ust_rst_ete_mult_retire_sys_ip               ),
    .ust_en_sys_op         ( ust_en_ete_mult_retire_sys_op                ),
    .ust_us_msg_data_ip    ( ust_ete_mult_retire_us_msg_data_w            ),
    .ust_us_msg_event_ip   ( ust_ete_mult_retire_us_msg_event_w           ),
    .ust_us_msg_ready_op   ( ust_ete_mult_retire_us_msg_ready_w           ),
    .ust_us_msg_valid_ip   ( ust_ete_mult_retire_us_msg_valid_w           ),
    .ust_ds_msg_data_op    ( ust_ete_mult_retire_ds_msg_data_w            ),
    .ust_ds_msg_event_op   ( ust_ete_mult_retire_ds_msg_event_w           ),
    .ust_ds_msg_ready_ip   ( ust_ete_mult_retire_ds_msg_ready_w           ),
    .ust_ds_msg_valid_op   ( ust_ete_mult_retire_ds_msg_valid_w           ),
    .ust_gpio_output_op    ( ust_ete_mult_retire_gpio_output_op           ),
    .ust_rv_halted_ip      ( ust_ete_mult_retire_rv_halted_ip             ),
    .ust_rv_stall_op       ( ust_ete_mult_retire_rv_stall_op              ),
    .ust_rv_i_retire_ip    ( ust_ete_mult_retire_rv_i_retire_ip           ),
    .ust_rv_i_lastsize_ip  ( ust_ete_mult_retire_rv_i_lastsize_ip         ),
    .ust_rv_i_type_ip      ( ust_ete_mult_retire_rv_i_type_ip             ),
    .ust_rv_i_sijump_ip    ( ust_ete_mult_retire_rv_i_sijump_ip           ),
    .ust_rv_i_uiret_ip     ( ust_ete_mult_retire_rv_i_uiret_ip            ),
    .ust_rv_i_address_ip   ( ust_ete_mult_retire_rv_i_address_ip          ),
    .ust_rv_i_context_ip   ( ust_ete_mult_retire_rv_i_context_ip          ),
    .ust_rv_i_ctype_ip     ( ust_ete_mult_retire_rv_i_ctype_ip            ),
    .ust_rv_i_ecause_ip    ( ust_ete_mult_retire_rv_i_ecause_ip           ),
    .ust_rv_i_tval_ip      ( ust_ete_mult_retire_rv_i_tval_ip             ),
    .ust_rv_i_privilege_ip ( ust_ete_mult_retire_rv_i_privilege_ip        ),
    .ust_rv_i_trigger_ip   ( ust_ete_mult_retire_rv_i_trigger_ip          ),
    .ust_rv_i_impdef_ip    ( ust_ete_mult_retire_rv_i_impdef_ip           ),
    .ust_rv_i_status_ip    ( ust_ete_mult_retire_rv_i_status_ip           ),
    .ust_rv_i_enabled_op   ( ust_ete_mult_retire_rv_i_enabled_op          ),
    .ust_lock_ip           ( 1'd0                                         ),
    .ust_locked_op         (                                              ),
    .ust_instance_id_ip    ( ust_ete_mult_retire_instance_id_ip           ),
    .ust_version_op        ( ust_ete_mult_retire_version_op               ),
    .ust_testmode_ip       ( ust_ete_mult_retire_testmode_ip              ),
    .ust_test_in_0_ip      ( {(ete_mult_retire_test_in_0_width_p){1'b0}}  ),
    .ust_test_out_0_op     (                                              )
  );

endmodule
